package reg_bus_pkg;
   typedef enum logic [7:0] {IDLE = 0,WTR_RRD=1,CWL_CL=2,RP_RTP=3,WR=4,
			     BL_RCD=5,RAS=6,FAW=7,ZQS=8,AREF=9,AREF_1=10,
			     AREF_2=11,RFC=12,RFC_1=13,DRV_IMP_RON_DATA=14,
			     DRV_IMP_RON_ADDR=15,DRV_IMP_RTT_DATA=16,DRV_SLEW=17,
			     MR0=18,MR0_1=19,MR1=20,MR1_1=21,MR2=22,
			     MR2_1=23,MR3=24,MR3_1=25,RG_REF_START_ADDR=26,
			     RG_REF_START_ADDR_1=27,RG_REF_END_ADDR=28,
			     RG_REF_END_ADDR_1=29,RG_REF_NUM_ROW_PER_REF=30,
			     RG_REF_EN_RASMIN=31,RG_REF_RP_RRD=32,
			     DRV_OCD_CAL_PU=33,DRV_OCD_CAL_PD=34,
			     DRV_OCD_CAL_DIS=35,DQS_OFFSET=36,DQS_OFFSET_1=37,
			     CLK_OFFSET=38,CLK_OFFSET_1=39,DISABLE_REF=40,
			     TREG_END=41,DRV_END=42,MODE_END=43,RG_REF_END=44,
			     RD_STATUS_MC=45,RD_STATUS_PHY_10=46,
			     RD_STATUS_PHY_11=47,RD_STATUS_PHY_12=48,
			     RD_STATUS_PHY_13=49,RD_STATUS_PHY_20=50,
			     RD_STATUS_PHY_21=51,RD_STATUS_PHY_22=52,
			     RD_STATUS_PHY_23=53,RD_STATUS_INIT_1=54,
			     RD_STATUS_INIT_2=55,BYPASS_BUS_RDY=56,
			     DRV_DLL_CAL_DIS=57,CONGEN_C3=58,
			     CONGEN_C4=59,CONGEN_C5=60,
			     CONGEN_C6=61,CONGEN_C7=62,CONGEN_C8=63,
			     CONGEN_C9=64,CONGEN_C10=65,CONGEN_R0=66,
			     CONGEN_R1=67,CONGEN_R2=68,CONGEN_R3=69,
			     CONGEN_R4=70,CONGEN_R5=71,CONGEN_R6=72,
			     CONGEN_R7=73,CONGEN_R8=74,CONGEN_R9=75,
			     CONGEN_R10=76,CONGEN_R11=77,CONGEN_R12=78,
			     CONGEN_R13=79,CONGEN_R14=80,CONGEN_R15=81,
			     CONGEN_B0=82,CONGEN_B1=83,CONGEN_B2=84,
			     CONGEN_XOR_SEL=85,CONGEN_END=86} REG_BUS_FRAMES;
endpackage: reg_bus_pkg
